library WORK;

package GENERICS is

    -- No constants

end package;
