library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

library WORK;
use WORK.TOP_LEVEL_CONSTANTS.ALL;

entity MODULE_ID is

end entity;

architecture RTL of MODULE_ID is
        
begin   
    

end architecture;