library WORK;

package MODULES is

    -- No constants

end package;
