library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.MATH_REAL.ALL;
use std.textio.all;

library WORK;

entity GENERIC_ROM IS

    generic (
        DATA_WIDTH        : natural := 8;
        ADDRESS_WIDTH     : natural := 8;
        ADDRESSABLE_WIDTH : natural := 7;
        INIT_FILE         : string  := "../data/mif/generic_rom_dummy.mif"
    );

    port (
        address     : in  std_logic_vector((ADDRESS_WIDTH - 1) downto 0);
        destination : out std_logic_vector((DATA_WIDTH - 1) downto 0) 
    );

end entity;

architecture RTL of GENERIC_ROM is

    type memory_block is array(0 TO (2**ADDRESSABLE_WIDTH - 1)) of std_logic_vector((DATA_WIDTH - 1) DOWNTO 0);

    impure function memory_init return memory_block is
        file     text_file : text open read_mode is INIT_FILE;
        variable text_line : line;
        variable content   : memory_block;
        variable index     : integer := 0;
        variable value     : bit_vector((DATA_WIDTH - 1) DOWNTO 0);
    begin
        while not endfile(text_file) loop
            readline(text_file, text_line);
            read(text_line, index);
            read(text_line, value);

            if index >= 0 and index < (2**ADDRESSABLE_WIDTH) then
                content(index) := To_StdLogicVector(value);
            end if;
        end loop;
        
        return content;
    end function;

    signal memory_ROM : memory_block := memory_init;

begin

    process(address)
        variable index : natural;
    begin
        index := to_integer(unsigned(address));
        if (index < (2**ADDRESSABLE_WIDTH - 1)) then
            destination <= memory_ROM(index);
        else
            destination <= (others => '0');
        end if;
    end process;

end architecture;
